library verilog;
use verilog.vl_types.all;
entity tb_stpm_full_sv_unit is
end tb_stpm_full_sv_unit;
