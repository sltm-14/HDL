library verilog;
use verilog.vl_types.all;
entity tb_mux_param is
end tb_mux_param;
