library verilog;
use verilog.vl_types.all;
entity ff_d_pkg is
end ff_d_pkg;
