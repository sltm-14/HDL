library verilog;
use verilog.vl_types.all;
entity mux_pkg is
end mux_pkg;
