library verilog;
use verilog.vl_types.all;
entity TB_bcd_7seg is
end TB_bcd_7seg;
