library verilog;
use verilog.vl_types.all;
entity tb2_ALU is
end tb2_ALU;
