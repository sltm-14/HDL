library verilog;
use verilog.vl_types.all;
entity tb_bin_to_dec is
end tb_bin_to_dec;
