`timescale 1ns / 1ps

module pwm #(parameter TOTAL_BITS = 8, POL = 1)
(
    input                       iClk,
    input                       iCE,
    input                       iRst,
    input   [(TOTAL_BITS-1):0]  ivDutyCycle,

    output                      oPWM,
    output                      oCycleStart
);
//////////////////////////////////////////////////////////////////////////////////
// Includes
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Defines
//////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////
// Internal Signals
//////////////////////////////////////////////////////////////////////////////////
//!
reg                         rPWM_d;
reg                         rPWM_q;
//!
reg     [(TOTAL_BITS-1):0]  rvCnt_d;
reg     [(TOTAL_BITS-1):0]  rvCnt_q;
//!
reg                         rCycleStart_d;
reg                         rCycleStart_q;
//////////////////////////////////////////////////////////////////////////////////
// Continous assigment
//////////////////////////////////////////////////////////////////////////////////
assign  oPWM        =   rPWM_q;
assign  oCycleStart =   rCycleStart_q;
//////////////////////////////////////////////////////////////////////////////////
// Sequential Section
//////////////////////////////////////////////////////////////////////////////////
always @(posedge iClk or posedge iRst)
begin
    if(iRst)
    begin
        rPWM_q          <=  ~POL;
        rvCnt_q         <=  {TOTAL_BITS{1'b0}};
        rCycleStart_q   <=  1'b0;
    end
    else
    begin
        rPWM_q          <=  rPWM_d;
        rCycleStart_q   <=  rCycleStart_d;
        if(iCE)begin
            rvCnt_q     <=  rvCnt_d;
        end
        else begin
            rvCnt_q     <=  rvCnt_q;
        end
    end
end
//////////////////////////////////////////////////////////////////////////////////
// Combinational Section
//////////////////////////////////////////////////////////////////////////////////
always @*
begin
    rvCnt_d         =   rvCnt_q + 1'b1  ;
    rPWM_d          =   (rvCnt_q < ivDutyCycle) ? ~POL : POL;
    rCycleStart_d   =   ~|rvCnt_q;
end
//////////////////////////////////////////////////////////////////////////////////
//Instances
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
endmodule
