library verilog;
use verilog.vl_types.all;
entity tb_ff_d is
end tb_ff_d;
