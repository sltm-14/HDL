library verilog;
use verilog.vl_types.all;
entity tb_pipo is
end tb_pipo;
