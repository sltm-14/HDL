library verilog;
use verilog.vl_types.all;
entity tb_dec_to_bin is
end tb_dec_to_bin;
