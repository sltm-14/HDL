`ifndef FF_D_PKG
    `define FF_D_PKG

    package ff_d_pkg;

        localparam DW = 4;

        typedef logic [DW-1:0] t_dw;

    endpackage

`endif
