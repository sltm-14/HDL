library verilog;
use verilog.vl_types.all;
entity tb_stpm_full is
end tb_stpm_full;
